[aimspice]
[description]
163
Double alternating rectifier
D1 a b DiodaSi
R b 0 100
D2 0 a DiodaSi
D3 0 c DiodaSi
D4 c b DiodaSi
.Model DiodaSi D tt = 1e-9
Vin a c sin(0 10 1k 0 0)



[tran]
1e-9
6e-3
0
0.00001
0
[ana]
4 3
0
1 1
1 1 -2 10
3
v(a)
v(b)
v(c)
0
1 1
1 1 -2 10
1
v(b)
0
1 1
1 1 -2 10
2
v(a)
v(c)
[end]
