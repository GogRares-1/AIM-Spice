[aimspice]
[description]
306
Reaction regulator with no error amplifier 
D1 a b DiodaSi
R outr 0 100
C b 0 1m
D2 0 a DiodaSi
D3 0 c DiodaSi
D4 c b DiodaSi
D5 0 z Zener
R1 b z 220
Q1 b z outr tranzistor

.Model DiodaSi D tt = 1e-9
.Model Zener D bv=5.6
.Model tranzistor NPN tr=1e-9 tf=1e-9
Vin a c DC 5 sin(0 10 50 0 0)

[tran]
1e-9
60e-3
X
X
0
[ana]
4 1
0
1 1
1 1 -3.41661E-22 5
1
v(outr)
[end]
