[aimspice]
[description]
125
Mono alternating rectifier ( Half waves )
D1 a b DiodaSi
.Model DiodaSi D tt = 1e-9
RL b 0 100
Vin a 0 sin(0 10 1k 0 0)

[tran]
1e-9
6e-3
0
0.00001
0
[ana]
4 1
0
1 1
1 1 -10 10
2
v(a)
v(b)
[end]
