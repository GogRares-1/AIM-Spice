[aimspice]
[description]
251
transmission gate
Vdd dd 0 DC 5
Vss ss 0 DC 0
Vap ap 0 DC 0
Van an 0 DC 5
Vin a 0 DC 0 pulse(0 5 0 1e-10 1e-10 1e-6 2e-6)
!
mp a an out dd cmos2 l=10u w=1u
mn a ap out ss cmos l=10u w=1u
!
.model cmos nmos vto=1.5
.model cmos2 pmos vto=-1.5
[dc]
1
Vin
0
5
0.1
[tran]
1e-9
6e-6
X
X
0
[ana]
1 2
0
1 1
1 1 0 5
1
v(out)
0
1 1
1 1 0 5
1
vin
[end]
