[aimspice]
[description]
220
Parametric regulator with Zener diode
D1 a b DiodaSi
R b 0 100
C b 0 1m
D2 0 a DiodaSi
D3 0 c DiodaSi
D4 c b DiodaSi
D5 0 b Zener
.Model DiodaSi D tt = 1e-9
.Model Zener D bv=6.8
Vin a c DC 5 sin(0 10 50 0 0)

[tran]
1e-9
60e-3
X
X
0
[ana]
4 1
0
1 1
1 1 -3.44663E-29 8
1
v(b)
[end]
