[aimspice]
[description]
191
NMOS
!
.model t1 nmos vto=1.5
.model t2 nmos vto=2.5
!
VGG g 0 7.5
VDD d 0 5
VIN in 0 DC pulse(0 5 0 1e-10 1e-10 1e-9 2e-9)
!
m1 OUT in 0 0 t1 l=1u W=1u
m2 d g OUT OUT t2 l=10u W=1u
[dc]
1
VIN
0
5
0.1
[tran]
1e-10
6e-9
X
X
0
[ana]
1 0
[end]
